.title KiCad schematic
R2 out1 Net-_R2-Pad2_ 10k
v1 Net-_R2-Pad2_ GND DC
v2 in GND sine
U2 out1 plot_v1
X1 unconnected-_X1-Pad1_ out1 Net-_R2-Pad2_ in GND unconnected-_X1-Pad6_ unconnected-_X1-Pad7_ unconnected-_X1-Pad8_ unconnected-_X1-Pad9_ unconnected-_X1-Pad10_ unconnected-_X1-Pad11_ GND unconnected-_X1-Pad13_ unconnected-_X1-Pad14_ BA10339F
.end
