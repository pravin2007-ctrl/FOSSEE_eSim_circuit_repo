.title KiCad schematic
U1 unconnected-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ unconnected-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ unconnected-_U1-Pad14_ PORT
U13 Net-_U13-Pad1_ Net-_U13-Pad2_ d_inverter
U12 Net-_U12-Pad1_ Net-_U12-Pad2_ d_inverter
U11 Net-_U11-Pad1_ Net-_U11-Pad2_ d_inverter
U4 Net-_U1-Pad5_ Net-_U10-Pad1_ d_inverter
U3 Net-_U1-Pad4_ Net-_U3-Pad2_ d_inverter
U7 Net-_U1-Pad9_ Net-_U13-Pad1_ d_inverter
U6 Net-_U1-Pad10_ Net-_U12-Pad1_ d_inverter
U5 Net-_U1-Pad11_ Net-_U11-Pad1_ d_inverter
U2 Net-_U1-Pad3_ Net-_U2-Pad2_ d_inverter
U9 Net-_U3-Pad2_ Net-_U14-Pad2_ d_inverter
U8 Net-_U2-Pad2_ Net-_U14-Pad1_ d_inverter
U10 Net-_U10-Pad1_ Net-_U10-Pad2_ d_inverter
U14 Net-_U14-Pad1_ Net-_U14-Pad2_ Net-_U14-Pad3_ d_and
U17 Net-_U1-Pad2_ Net-_U17-Pad2_ d_inverter
U21 Net-_U17-Pad2_ Net-_U21-Pad2_ d_inverter
U16 Net-_U1-Pad13_ Net-_U16-Pad2_ d_inverter
U20 Net-_U16-Pad2_ Net-_U20-Pad2_ d_inverter
U18 Net-_U14-Pad3_ Net-_U10-Pad2_ Net-_U18-Pad3_ d_and
U15 Net-_U11-Pad2_ Net-_U12-Pad2_ Net-_U15-Pad3_ d_and
U19 Net-_U15-Pad3_ Net-_U13-Pad2_ Net-_U19-Pad3_ d_and
U26 Net-_U24-Pad2_ Net-_U1-Pad6_ d_inverter
U25 Net-_U23-Pad2_ Net-_U1-Pad8_ d_inverter
U23 Net-_U22-Pad6_ Net-_U23-Pad2_ d_inverter
U24 Net-_U22-Pad7_ Net-_U24-Pad2_ d_inverter
U22 Net-_U18-Pad3_ Net-_U19-Pad3_ Net-_U1-Pad12_ Net-_U20-Pad2_ Net-_U21-Pad2_ Net-_U22-Pad6_ Net-_U22-Pad7_ d_jkff
.end
